module ASYN_FIFO (

);





endmodule