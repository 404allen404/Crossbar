module ID_Decoder (


);



endmodule
