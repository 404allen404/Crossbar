module RPTR_EMPTY ();



endmodule