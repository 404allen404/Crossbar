module AXI_M_IF (


);


endmodule